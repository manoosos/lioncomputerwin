version https://git-lfs.github.com/spec/v1
oid sha256:e7e43462353a5ee296d1b2114d20ea9f89c7c47aa59ac6c100313ec8718524fa
size 33554944
